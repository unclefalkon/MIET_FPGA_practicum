module fsm(
    input clk100_i,
    input rstn_o
);

endmodule