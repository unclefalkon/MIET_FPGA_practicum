module stopwatch(
    input clk100_i,
    input rstn_i,
    input start_stop_i,
    output [6:0] hex0_o,
    output [6:0] hex1_o,
    output [6:0] hex2_o,
    output [6:0] hex3_o
);

endmodule