module fsm_with_fifo(
    input clk100_i,
    input rstn_i,
    input [7:0] data_i,
    input we_i,
    output full_o,
    output transmit_lane_o
);

endmodule