module ps2_ctrl(
    input clk100_i,
    input rstn_i,
    input ps2_clk_i,
    input ps2_dat_i,

    output reg valid_data_o,
    output [7:0] data_o
);

endmodule