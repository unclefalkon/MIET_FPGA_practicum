module stopwatch(
    input start_stop,
    input reset,
    input clk,
    output [6:0] HEX0,
    output [6:0] HEX1,
    output [6:0] HEX2,
    output [6:0] HEX3
);

endmodule